// This file is where you'll define the testbench for your simple ALU 
// for project 1. Refer to the project one document for instructions 
// and guidance.

`timescale 10ms/1ms

module ALU_testbench();

// Instantiate your ALU and implement your testbench here

endmodule