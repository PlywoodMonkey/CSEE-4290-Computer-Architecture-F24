
// This file is where you'll define your simple ALU for project 1.
// Refer to the project one document for instructions and guidance.

module ALU
(
    // Input/Output definitions here
);

// Implementation here

endmodule